library verilog;
use verilog.vl_types.all;
entity keyscan_vlg_tst is
end keyscan_vlg_tst;
